//UVM sequence items