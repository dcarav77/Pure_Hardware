//UVM environment